library verilog;
use verilog.vl_types.all;
entity NLC_testbench_stud is
end NLC_testbench_stud;
