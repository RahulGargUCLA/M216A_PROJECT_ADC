library verilog;
use verilog.vl_types.all;
entity NLC_6th_order_16ch_testbench is
end NLC_6th_order_16ch_testbench;
